../ex4.5/ex405.sv